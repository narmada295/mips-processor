module andm(inA, inB, out);
    input inA, inB;
    output out;
    
    and and_gate(out, inA, inB);
endmodule
